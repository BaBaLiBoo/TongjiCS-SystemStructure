`timescale 1ns / 1ps

module Register_IF_ID (
    input  wire        clk_i,
    input  wire        rst_i,
    input  wire        stall_i,  // ͣ���ź�
    input  wire        branch_i, // ��֧ˢ���ź�
    input  wire [31:0] npc_i,
    input  wire [31:0] instruction_i,
    
    output reg  [31:0] npc_o,
    output reg  [31:0] instruction_o
);

    always @(posedge clk_i or posedge rst_i) begin
        if (rst_i) begin
            npc_o <= 32'b0;
            instruction_o <= 32'b0;
        end 
        else if (stall_i) begin
            // ͣ��
            if (branch_i) begin
                npc_o <= 32'b0;
                instruction_o <= 32'b0;
            end
            else begin
                // ���ֲ���
                npc_o <= npc_o;
                instruction_o <= instruction_o;
            end
        end 
        else if (branch_i) begin
            // ��֧ˢ��
            npc_o <= 32'b0;
            instruction_o <= 32'b0; // ע�� nop
        end
        else begin
            // ��������
            npc_o <= npc_i;
            instruction_o <= instruction_i;
        end
    end

endmodule