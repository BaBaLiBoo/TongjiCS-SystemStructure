`define STATUS          12
`define CAUSE           13
`define EPC             14
`define CAUSE_SYSCALL   5'b01000
`define CAUSE_BREAK     5'b01001
`define CAUSE_TEQ       5'b01101

`define OPC_ADDI        6'b001000
`define OPC_ADDIU       6'b001001
`define OPC_ANDI        6'b001100
`define OPC_ORI         6'b001101
`define OPC_SLTIU       6'b001011
`define OPC_LUI         6'b001111
`define OPC_XORI        6'b001110
`define OPC_SLTI        6'b001010
`define OPC_ADDU        6'b000000
`define OPC_AND         6'b000000
`define OPC_BEQ         6'b000100
`define OPC_BNE         6'b000101
`define OPC_JR          6'b000000
`define OPC_LW          6'b100011
`define OPC_XOR         6'b000000
`define OPC_NOR         6'b000000
`define OPC_OR          6'b000000
`define OPC_SLL         6'b000000
`define OPC_SLLV        6'b000000
`define OPC_SLTU        6'b000000
`define OPC_SRA         6'b000000
`define OPC_SRL         6'b000000
`define OPC_SUBU        6'b000000
`define OPC_SW          6'b101011
`define OPC_ADD         6'b000000
`define OPC_SUB         6'b000000
`define OPC_SLT         6'b000000
`define OPC_SRLV        6'b000000
`define OPC_SRAV        6'b000000
`define OPC_CLZ         6'b011100
`define OPC_DIVU        6'b000000
`define OPC_ERET        6'b010000
`define OPC_LHU         6'b100101
`define OPC_SB          6'b101000
`define OPC_SH          6'b101001
`define OPC_LH          6'b100001
`define OPC_MFHI        6'b000000
`define OPC_MFLO        6'b000000
`define OPC_MTHI        6'b000000
`define OPC_MTLO        6'b000000
`define OPC_MUL         6'b011100
`define OPC_MULTU       6'b000000
`define OPC_SYSCALL     6'b000000
`define OPC_TEQ         6'b000000
`define OPC_BGEZ        6'b000001
`define OPC_BREAK       6'b000000
`define OPC_DIV         6'b000000
`define OPC_J           6'b000010
`define OPC_JAL         6'b000011
`define OPC_JALR        6'b000000
`define OPC_LB          6'b100000
`define OPC_LBU         6'b100100

`define FNC_ADDU        6'b100001
`define FNC_AND         6'b100100
`define FNC_JR          6'b001000
`define FNC_XOR         6'b100110
`define FNC_NOR         6'b100111
`define FNC_OR          6'b100101
`define FNC_SLL         6'b000000
`define FNC_SLLV        6'b000100
`define FNC_SLTU        6'b101011
`define FNC_SRA         6'b000011
`define FNC_SRL         6'b000010
`define FNC_SUBU        6'b100011
`define FNC_ADD         6'b100000
`define FNC_SUB         6'b100010
`define FNC_SLT         6'b101010
`define FNC_SRLV        6'b000110
`define FNC_SRAV        6'b000111
`define FNC_CLZ         6'b100000
`define FNC_DIVU        6'b011011
`define FNC_ERET        6'b011000
`define FNC_JALR        6'b001001
`define FNC_MFHI        6'b010000
`define FNC_MFLO        6'b010010
`define FNC_MTHI        6'b010001
`define FNC_MTLO        6'b010011
`define FNC_MUL         6'b000010
`define FNC_MULTU       6'b011001
`define FNC_SYSCALL     6'b001100
`define FNC_TEQ         6'b110100
`define FNC_BREAK       6'b001101
`define FNC_DIV         6'b011010
